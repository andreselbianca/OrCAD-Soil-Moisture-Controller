** Profile: "SCHEMATIC1-ParametricConvertor"  [ d:\an 2-etti\tehnici cad-proiecte orcad\proiectcad-PSpiceFiles\SCHEMATIC1\ParametricConvertor.sim ] 

** Creating circuit file "ParametricConvertor.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../blueled.lib" 
* From [PSPICE NETLIST] section of C:\Users\bianca\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5s 0 1m 
.STEP LIN PARAM r 600k 100k 100k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
